LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.STD_LOGIC_UNSIGNED.ALL;
LIBRARY displayNumber;
ENTITY part5 IS
	PORT(SW: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		  HEX0: OUT STD_LOGIC_VECTOR(0 TO 6);
		  HEX1: OUT STD_LOGIC_VECTOR(0 TO 6);
		  HEX2: OUT STD_LOGIC_VECTOR(0 TO 6);
		  HEX3: OUT STD_LOGIC_VECTOR(0 TO 6);
		  LEDR: OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
		  
END part5;


ARCHITECTURE Structure of part5 IS
	COMPONENT displayNumber IS
		PORT(s	:IN	STD_LOGIC_VECTOR(0 TO 3);
			  HEX	:OUT	STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;
	COMPONENT fulladder IS
		PORT(Cin: IN STD_LOGIC;
			A: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			O: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			Cout: OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT displayTwoNumbers IS
		PORT(L: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  C: IN STD_LOGIC;
		  HEX1: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		  HEX0: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
	END COMPONENT;
	SIGNAL display: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL TEMPC: STD_LOGIC;
BEGIN 
	stage0: LEDR<=SW;
	stage1: displayNumber PORT MAP(SW(7 DOWNTO 4),HEX3);
	stage2: displayNumber PORT MAP(SW(3 DOWNTO 0),HEX2);
	stage3: fulladder PORT MAP('0',SW(7 DOWNTO 4),SW(3 DOWNTO 0),display,TEMPC);
	stage4: displayTwoNumbers PORT MAP(display,TEMPC,HEX1,HEX0);
END Structure;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.STD_LOGIC_UNSIGNED.ALL;
ENTITY fulladder IS
	PORT(Cin: IN STD_LOGIC;
			A: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			O: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			Cout: OUT STD_LOGIC);
END fulladder;

ARCHITECTURE LogicFunction OF fulladder IS
	SIGNAL Z,TEMPC,Q,T,V:STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN 
	TEMPC<="0000" & Cin;
	Q<= ('0'&A)+('0'&B);
	T <= TEMPC +Q;
	PROCESS(T
	)
	BEGIN
		IF T>"1001" THEN
			Z<= "01010";
			Cout <= '1';
		ELSE
			Z<="00000";
			Cout<='0';
		END IF;
	END PROCESS;
	V<= T-Z;
	O<=V(3 DOWNTO 0);
END LogicFunction;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.STD_LOGIC_UNSIGNED.ALL;

ENTITY displayTwoNumbers IS
	PORT(L: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  C: IN STD_LOGIC;
		  HEX1: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		  HEX0: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END displayTwoNumbers;

ARCHITECTURE LogicFunction OF displayTwoNumbers IS
	SIGNAL T,N: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL H: STD_LOGIC;
BEGIN
	N<=L;
	PROCESS(C)
	BEGIN
	IF C='0' THEN
		HEX1<="0000001";
	ELSE      
		HEX1<="1001111";
	END IF;
	END PROCESS;
	PROCESS(T)
	BEGIN
	CASE N IS 
				WHEN "0000" => HEX0<="0000001";
				WHEN "0001" => HEX0<="1001111";
				WHEN "0010" => HEX0<="0010010";
				WHEN "0011" => HEX0<="0000110";
				WHEN "0100" => HEX0<="1001100";
				WHEN "0101" => HEX0<="0100100";
				WHEN "0110" => HEX0<="0100000";
				WHEN "0111" => HEX0<="0001111";
				WHEN "1000" => HEX0<="0000000";
				WHEN "1001" => HEX0<="0000100";
				WHEN OTHERS => HEX0<="-------";
	END CASE;
	END PROCESS;	
		
	  
		
		




END LogicFunction;




		
