LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY bit4_counter IS
	PORT(En,CLK,CLR: IN STD_LOGIC;
					Q1,Q2,Q3,Q4: OUT STD_LOGIC:='0');
END bit4_counter;

ARCHITECTURE structure OF bit4_counter IS
	COMPONENT T_FF
		PORT(T,CLK,CLR : IN STD_LOGIC;
					Q : OUT STD_LOGIC);
	END COMPONENT;	
	SIGNAL C1,C2,C3: STD_LOGIC;
	SIGNAL TMP: STD_LOGIC_VECTOR(1 TO 4):="0000";
BEGIN
	STAGE1: T_FF PORT MAP(EN,CLK,CLR,TMP(1));
	STAGE1_2: C1 <= EN AND TMP(1);
	STAGE2: T_FF PORT MAP(C1,CLK,CLR,TMP(2));
	STAGE2_2: C2 <= TMP(2) AND C1;
	STAGE3: T_FF PORT MAP(C2,CLK,CLR,TMP(3));
	STAGE3_2: C3 <= TMP(3) AND C2;
	STAGE4: T_FF PORT MAP(C3,CLK,CLR,TMP(4));
	STAGE5: Q4 <= TMP(4);
	STAGE6: Q3 <= TMP(3);
	STAGE7: Q2 <= TMP(2);
	STAGE8: Q1 <= TMP(1);
END structure;