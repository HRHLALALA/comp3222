LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY displayNumber;
LIBRARY adder4;
LIBRARY Comparator;
LIBRARY part2;

ENTITY part4 IS
	PORT(SW: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		  LEDR: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		  HEX0: OUT STD_LOGIC_VECTOR(0 TO 6);
		  HEX1: OUT STD_LOGIC_VECTOR(0 TO 6);
		  HEX2: OUT STD_LOGIC_VECTOR(0 TO 6);
		  HEX3: OUT STD_LOGIC_VECTOR(0 TO 6);
		  LEDG: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END part4;

ARCHITECTURE STRUCTURE OF part4 IS
	COMPONENT displayNumber IS
		PORT(s	:IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
			  HEX	:OUT	STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;
	COMPONENT Comparator IS
		PORT (X:	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Z: OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT adder4 IS
		PORT(Cin	:IN STD_LOGIC;
			X	:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Y	:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			S	:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			Cout: OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT part2 IS
		PORT ( SW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
					C: IN STD_LOGIC;
				HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6);
				HEX1 : OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;
	SIGNAL TEMP1,TEMP2,CARRY: STD_LOGIC;
	SIGNAL RESULT: STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	init1: LEDR<=SW;
	init2: displayNumber PORT MAP(SW(7 DOWNTO 4),HEX3);
	init3: displayNumber PORT MAP(SW(3 DOWNTO 0),HEX2);
	init4: Comparator PORT MAP(SW(7 DOWNTO 4),TEMP1);
	init5: Comparator PORT MAP(SW(3 DOWNTO 0),TEMP2);
	init6: LEDG(7)<= TEMP1 OR TEMP2;
	stage0: adder4 PORT MAP('0',SW(3 DOWNTO 0),SW(7 DOWNTO 4),RESULT,CARRY);
	stage1: LEDG(3 DOWNTO 0)<=RESULT;
	stage2: LEDG(4)<= CARRY;
	stage3: part2 PORT MAP(RESULT,CARRY,HEX0,HEX1);
	
	



END STRUCTURE;
	