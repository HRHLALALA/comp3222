LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY part4 IS
	PORT(D,Clock: 	IN STD_LOGIC;
			Qa,Qb,Qc: OUT STD_LOGIC;)
			
ARCHITECTURE 
			