LIBRARY ieee;
USE ieee. std_logic_1164.all;

ENTITY part1 IS
	PORT(En,CLK,CLR: IN STD_LOGIC;
			Q: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END part1;

ARCHITECTURE Structure OF part1 IS
	COMPONENT T_FF
		PORT(T,CLK,CLR : IN STD_LOGIC;
					Q : OUT STD_LOGIC);
	END COMPONENT;	 
	SIGNAL TMP: STD_LOGIC_VECTOR(8 DOWNTO 1);
	SIGNAL C1,C2,C3,C4,C5,C6,C7: STD_LOGIC;
BEGIN
	STAGE1: T_FF PORT MAP(EN,CLK,CLR,TMP(1));
	STAGE1_2: C1 <= EN AND TMP(1);
	STAGE2: T_FF PORT MAP(C1,CLK,CLR,TMP(2));
	STAGE2_2: C2 <= TMP(2) AND C1;
	STAGE3: T_FF PORT MAP(C2,CLK,CLR,TMP(3));
	STAGE3_2: C3 <= TMP(3) AND C2;
	STAGE4: T_FF PORT MAP(C3,CLK,CLR,TMP(4));
	STAGE4_2: C4 <= TMP(4) AND C3;
	STAGE5: T_FF PORT MAP(C4,CLK,CLR,TMP(5));
	STAGE5_2: C5 <= TMP(5) AND C4;
	STAGE6: T_FF PORT MAP(C5,CLK,CLR,TMP(6));
	STAGE6_2: C6 <= TMP(6) AND C5;
	STAGE7: T_FF PORT MAP(C6,CLK,CLR,TMP(7));
	STAGE7_2: C7 <= TMP(7) AND C6;
	STAGE8: T_FF PORT MAP(C7,CLK,CLR,TMP(8));
	STAGE9: Q<=TMP;
END Structure;
	
		