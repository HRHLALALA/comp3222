LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY D_FF IS
	PORT(D,CLOCK:IN STD_LOGIC;
			Q		:OUT STD_LOGIC);
END D_FF;

ARCHITECTURE Behavior OF D_FF IS
BEGIN
	PROCESS(CLOCK)
	BEGIN
		IF CLOCK'EVENT AND CLOCK ='1' THEN
			Q <= D;
		END IF;
	END PROCESS;
	
END Behavior;