library verilog;
use verilog.vl_types.all;
entity search_vlg_vec_tst is
end search_vlg_vec_tst;
