library verilog;
use verilog.vl_types.all;
entity bit4_counter_vlg_vec_tst is
end bit4_counter_vlg_vec_tst;
